package core0_pkg;


endpackage
