module alu (
    input logic [ 3:0] alu_ctrl,
    input logic [31:0] src1,
    input logic [31:0] src2,

    output logic [31:0] alu_res,
    output logic zero,
    output logic last_bit
);
  wire [4:0] shamt = src2[4:0];

  always_comb begin
    case (alu_ctrl)
      // ADD
      4'b0000: alu_res = src1 + src2;
      // AND
      4'b0010: alu_res = src1 & src2;
      // OR
      4'b0011: alu_res = src1 | src2;
      // SUB
      4'b0001: alu_res = src1 + (~src2 + 1'b1);  // -a = (~a+1) 2's complement
      // SLT
      4'b0101: alu_res = {31'b0, $signed(src1) < $signed(src2)};
      // SLTU
      4'b0111: alu_res = {31'b0, src1 < src2};
      // XOR
      4'b1000: alu_res = src1 ^ src2;
      // SLL
      4'b0100: alu_res = src1 << shamt;
      // SRL
      4'b0110: alu_res = src1 >> shamt;
      // SRA
      4'b1001: alu_res = $signed(src1) >>> shamt;
      default: alu_res = 32'd0;
    endcase
  end

  assign zero = alu_res == 32'd0;
  assign last_bit = alu_res[0];
endmodule
